`define ANALOG_BIT_SIZE 4
`define WAVE_LENGTH 4096
